`timescale 1ns/100ps

module through_module(
    input [15:0] i_input,
    output logic [15:0] o_output
);

initial begin 

end 


    assign o_output = i_input;

endmodule