`timescale 1ns/1ps

module axi_stream_source(
    input aclk;
    output tvalid;
    input tready;
    output [7:0] tdata;
);

endmodule